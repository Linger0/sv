module min_delay (
  input  a,
  input  b,
  output c
);
  assign c = a + b;
endmodule
